/*
 * Module Name: mod_sub
 * Author(s):
 * Target: FIPS 203 (ML-KEM / Kyber)
 *
 * Description:
 */

module mod_sub(

);

endmodule
